     
 LS Library                                   �          A                            
 LS Library                                  �        B                            
 LS Library                                  �        C                            
 LS Library          $                        �        D                            =
 LS Library       $ $                        �         ��         ��    �        ��      =
 LS Library       $                         �         �~         �~    �        ��      =
 LS Library       $                         �         |r         |r    �      	  ��      =
 LS Library       $                          �         �l         �l    �   
     ��      D
 LS Library       0                         �         �         �    �         �j         �j    �         �          �     �              ��      	 D
 LS Library       0                         �         i         i    �         Z�         Z�    �   	      "�         "�    �              ��      
 D
 LS Library       0                         �         ^7         ^7    �         ��         ��    �   
      B9         B9    �              ��       D
 LS Library       0 $                        �         ��         ��    �          ��         ��    �         B�         B�    �              ��       M
 LS Library       8                          �         b�         b�    �         �         �    �   -   .   /  ��(       M
 LS Library       8  
                       �   	      ^         ^    �         Ɛ         Ɛ    �   0   1   2  ��(       M
 LS Library       @                         �         XU         XU    �          �          �    �   3   4   5  ��(       
 LS Library         F                         �   <     g                                                                 	   
                   
                     	                
    	                  	  	       
  
                                              . .        )  ' (          '  $        	   
          !  	 "  !   " #  #      $   ! %  %   # &  &       $  (   
 )  ) *  *   & +  +   ( ,    6 ! ,  " 6 0 # 7  $ 7 1 %  8 & 8 - ' 9  ( 9 . ) 2 : * : 3 + ; / , ; 4 - 5 < = =                                           %           $ %           ) %           $            )            $            	 )           
 $             )            0            0           0           5        %    0   	         0   	        0   	        5   	     #  	  0   
         0   
        0   
    
    5   
        
  0 %           0 &      !    0 '           5 &       '    !           !          , %     	    ,     	 
     /          ! /          " .         # .          $ !          % /         & .          ' -         ( -          ) #           * # '         + . %        , - &     !   - 8 !       &   . 8 #      (   / = "       +   0 8        "  
 1 8       $  	 2 =        )   3 @        *   4 @       ,   5 E        -   6 5       "  
 7 5     # $  	 8 5 !    % &   9 5 #    ' (   : =     ) *   ; =     + ,   < F        -         2   7-SEGMENT DISPLAY (g)        A      B     C     D     g                      P xd       �An                                                        