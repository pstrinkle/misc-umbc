     
 LS Library 	      $         &          &     �         ��         ��    �         J�         J�    �         ��         ��    �         ��         ��    �         V�         V�    �         �         �    �         N�         N�    �         �u         �u    �   	      l         l    �   
      �         �    �         �<         �<    �         ��         ��    �          V          V    �         r�         r�    �         �         �    �         �         �    �         ��         ��    �         ��         ��    �         ��         ��    �         �"         �"    �         Đ         Đ    �         �P         �P    �         r�         r�    �         ҥ         ҥ    �         &�         &�    �                 �� ��C 8-BITFA2.CKT C:\CIRCUITS\8-BITFA2.CKT 8-BITFA2.CKTA � �V�    B � �V�   C-in  �V�   Sum   �V�    C-out �V�   ����������������������������������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
  ���� 
 LS Library	                �         �    �         �m         �m    �         �N         �N    �          �          �    �         �         �    �   	      2�         2�    �   
      |�         |�    �         �         �    �                      �         R�         R�    �         v         v    �         �5         �5    �         N          N     �         ��         ��    �                �� H��C 4-BITFA2.CKT C:\CIRCUITS\4-BITFA2.CKT 4-BITFA2.CKTA � �V�    B � �V�   C-in  �V�   Sum   �V�    C-out �V�   ����������������������������  �� �� �� �� �� �� �� �� ��
 �� �� �� �� ��  ���� 
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ���� `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                            ��     ��        ��       ��       ��       ��       ��       ��       ��           ��  	          
     ��                  ��                 ��        ��       ��   
 LS Library	               .P         .P    �         �         �    �         �          �     �         ƚ         ƚ    �         r         r    �                      �         @�         @�    �         �         �    �         jv         jv    �         �o         �o    �         b�         b�    �         �p         �p    �         ��         ��    �         �         �    �         	   
    �� H��C 4-BITFA2.CKT C:\CIRCUITS\4-BITFA2.CKT 4-BITFA2.CKTA out �V�    B out �V�   C-in  �V�   Sum   �V�    C-out �V�   ����������������������������  �� �� �� �� �� �� �� �� ��
 �� �� �� �� ��  ���� 
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ���� `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                            ��     ��        ��       ��       ��       ��       ��       ��       ��           ��  	          
     ��                  ��                 ��        ��       ��   `
 LS Library               ��         ��    �         ^�         ^�    �         b�         b�    �         {         {    �         n�         n�    �         �         �    �         ΐ         ΐ    �         ~�         ~�    �          .�         .�    �         ރ         ރ    �         �         �    �         ��         ��    �         �v         �v    �         �r         �r    �         Nn         Nn    �         ��         ��    �           ��                                                `
 LS Library              ^�         ^�    �   	      �>         �>    �   
      8�         8�    �         �         �    �         v.         v.    �         ��         ��    �         t�         t�    �         �         �    �         f         f    �   	      �         �    �   
      ��         ��    �         f         f    �                      �         V&         V&    �         $         $    �         �#         �#    �          ��                                               �� `
 LS Library       ,        �7         �7    �         :5         :5    �         �4         �4    �         ><         ><    �         �9         �9    �         �9         �9    �         @         @    �         �?         �?    �         ��         ��    �         T�         T�    �         ��         ��    �         `�         `�    �         V         V    �         *1         *1    �         �0         �0    �         �-         �-    �          !  ��                                               ����     ��         ��       ��       ��       ��        ��       ��       ��       ��     	  �� 	    
  �� 
      ��       ��       ��       ��       ��          ��        ��        ��       ��       ��                ��       ��       ��       ��       ��  ���� `
 LS Library       8 % #      T�         T�    �   $      T�         T�    �   %      ��         ��    �   &      ��         ��    �   #      
�         
�    �   $      x�         x�    �   %      �         �    �   &      T�         T�    �                 ��                                             
 LS Library                                   �         �         �    �         ��         ��    �         B�         B�    �         ��         ��    �         F�         F�    �         ��         ��    �         ��         ��    �   	    A                            
 LS Library                                  �   
     C-in                         
 LS Library                                  �         "         "    �         �9         �9    �         �=         �=    �         @A         @A    �          E          E    �          �         �    �   !      F         F    �   l    B                            
 LS Library         0        Z�         Z�    �         v�         v�    �         &�         &�    �         ��         ��    �         ��         ��    �         6�         6�    �         ��         ��    �         �p         �p    �        Sum                           
 LS Library         0        d�         d�    �        C-out                        	 `
 LS Library      / #       �w         �w    �         ή         ή    �         v         v    �         ��         ��    �         T�         T�    �         �         �    �         ��         ��    �         p�         p�    �   $  #  "  !      ��
                                            
 `
 LS Library      / '        �          �    �         ��         ��    �         ��         ��    �         0�         0�    �         ��         ��    �         ��         ��    �         ��         ��    �         ��         ��    �   )  (  '  &  %   ��
                                             
 LS Library	  	     2 !                        �         n;         n;    �         ;         ;    �         �:         �:    �         ~:         ~:    �         .:         .:    �         �9         �9    �         �9         �9    �   "      >9         >9    �   #     N �8        N �8    �   $      �8         �8    �   %      N8         N8    �   &      �7         �7    �   '      �7         �7    �   $   #   "   !   )   (   '   &   /           *  ��1  
 LS Library         A  (      ��         ��    �   )      ��         ��    �   *      �p         �p    �   +      ��         ��    �   #      ^�         ^�    �   $      �         �    �   %      ��         ��    �   &      n�         n�    �   8   	  Sum2                          
 LS Library         = ( '      ��         ��    �   9     Cout                          `
 LS Library       >  (      ��         ��    �   )      X�         X�    �   *      �         �    �   +      >�         >�    �   #      ��         ��    �   $      ��         ��    �   %      N�         N�    �   &      ��         ��    �   (      ��         ��    �   )      6�         6�    �   *      ��         ��    �   +      ��         ��    �   #      F�         F�    �   $      ��         ��    �   %      ��         ��    �   &      V�         V�    �   <   ;   8  ��                                               �� `
 LS Library       * $ (      ��         ��    �   )      h�         h�    �   *      �         �    �   +      Ȣ         Ȣ    �   (      x�         x�    �   )      (�         (�    �   *      ء         ء    �   +      ��         ��    �   D   C   B   A   @  ��                                             `
 LS Library      ! &       8�         8�    �   	      �         �    �   
      ��         ��    �         H�         H�    �         &�         &�    �   	      ֙         ֙    �   
      ��         ��    �         6�         6�    �   I  H  G  F  E   ��
                                             `
 LS Library      ! "        �         �    �         ��         ��    �         F�         F�    �         ��         ��    �          D�         D�    �         ��         ��    �         ��         ��    �         T�         T�    �   N  M  L  K  J   ��
                                             `
 LS Library       &       �         �    �   	      ��         ��    �   
      �         �    �         ��         ��    �         b�         b�    �         �         �    �                      �         r�         r�    �         "�         "�    �   	      p�         p�    �   
       �          �    �         �         �    �         �         �    �         0         0    �         �~         �~    �         �~         �~    �   Q  P  =   ��                                                `
 LS Library       "        @~         @~    �         �}         �}    �         �}         �}    �         P}         P}    �          }          }    �         �|         �|    �         `|         `|    �         |         |    �          �         �    �         ��         ��    �         f�         f�    �         �         �    �         ��         ��    �         v�         v�    �         &�         &�    �         ��         ��    �   T  S  R   ��                                               ������ 
 LS Library	  	     $                           �         n;         n;    �         ;         ;    �         �:         �:    �         ~:         ~:    �   	      .:         .:    �   
      �9         �9    �         �9         �9    �         >9         >9    �   (     N �8        N �8    �   )      �8         �8    �   *      N8         N8    �   +      �7         �7    �   "      �7         �7    �   N   M   L   K   I   H   G   F   ]   D  C  B  A  X  ��1  
 LS Library	               �         �    �         D�         D�    �         vc         vc    �         �b         �b    �         6b         6b    �         �a         �a    �          �`         �`    �   !      V`         V`    �         zB         zB    �         >;         >;    �   	      �:         �:    �   
      &C         &C    �         F@         F@    �         �?         �?    �         ?         ?    �         �_         �_    �         _         _    �      �   j  �� 6��C 8-BITXOR.CKT C:\CIRCUITS\8-BITXOR.CKT 8-BITXOR.CKTB � �V�    C-in  �V�   XOR'd �V�    ����������������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� 
 ���� ]
 LS Library                                  �         t�         t�    �   	      $�         $�    �           ��3        ]
 LS Library                                 �         ��         ��    �   
      ��         ��    �           ��3        ]
 LS Library                                 �         D�         D�    �         �         �    �      	   
  ��3        ]
 LS Library         %                        �         �y         �y    �         By         By    �           ��3        ]
 LS Library         +                        �         �k         �k    �         �k         �k    �           ��3        ]
 LS Library         0                        �         .^         .^    �         �]         �]    �           ��3        ]
 LS Library         6                        �         |P         |P    �         ,P         ,P    �           ��3       	 ]
 LS Library         ;                        �         �B         �B    �         zB         zB    �           ��3       
 `
 LS Library               8�         8�    �         �         �    �         �I         �I    �         �I         �I    �         >I         >I    �         �H         �H    �         �H         �H    �         NH         NH    �          �G         �G    �         �G         �G    �         ^G         ^G    �         G         G    �         �F         �F    �         nF         nF    �         F         F    �         �E         �E    �                  !      ��                                                                                 `
 LS Library       0  	      �D         �D    �   
      �B         �B    �         ~B         ~B    �         .B         .B    �         �A         �A    �         �A         �A    �         >A         >A    �         �@         �@    �   	      �@         �@    �   
      N@         N@    �         �?         �?    �         �?         �?    �         ^?         ^?    �         ?         ?    �         �>         �>    �         n>         n>    �   9   :   ;   <   =   >   ?   @   A  ��                                                                                ��     ��         ��        ��        ��        ��        ��        ��        ��  	     	 ��                       	   	      ��   
      ��        ��        ��        ��        ��        ��    	    ��  , ,                                                                                                                   	     	       
     
                                                                                                                                                                                                                                  !        "        #         $        %        &        '         (          )        *        +        N + ������            ��   ��������������������������������������������������������������( � R ) � � * � % + � � , � � - �   . � � / � � 0 � � 1 * 9 2 � / 3 � < 4 � � 5 �  6 � ; 7 @ � 8  � 9 � = : � � ; P � < Q E = S � > T J ? h � @ � � A � � B X � C � ] D f  E � � F    G g  H g h I  � J 	 f K 
 � L j � M l  � R   $         F            $        G   	 
       $            ,                    ,           ��������	         J           
  	       K            M          !       F D 8            0                   0           �� ,           	     I             ���������������� ; %       5  # $ % &  8 (           &  8 '           %  8 &           $  8 %             #   / #  	     -      ! 2 &  	          " 2 %  	          # 2 $  	          $ 2 #  	            % / '  
     *      & 2 *  
          ' 2 )  
          ( 2 (  
          ) 2 '  
           * 8 )      1  ' ��������/ 2 +      2  " ����������������8 A              ( ) * + # $ % & 9 = )       1  ' ��; >        6  # $ % & < >        3  ( ) * + =  &       9   	 
      ����@ - $       7  ( ) * + A * '           + B * &           * C * %           ) D * $             ( E ! &       <   	 
  F $ )            G $ (           
 H $ '           	 I $ &             J ! "       >       K $ %            L $ $            M $ #            N $ "               ��P  '      ;      Q  &       <   	 
  R  "       (           S  #      =      T  "       >       ������X * (      B  " ��������] $ *      C   ����������������f      J D           g "     H G   	 
      h "     H ?   	 
      ��j         L   	 
      ��l         M          ! ���������������������������������������������  "    8 (           �  &    : 9   	 
      �  *    @ C   �        A   � - '    * )      � - ,    , )      �   ,    , +      � - #    . -      � -     0 .      �       0 /      � .     4 3  ( ) * + � ;      6 5  # $ % & � . $    7 4  ( ) * + �      A E @   �   '    ; +      �   #    = /      �  	    I K E   � * +    B 2  " �      ? L :   	 
               Part 2       Part 1 
  ����   A     C-in     B     Sum     C-out  ��   Cout  	   Sum2                  	         P xd       �An                                                        