 
 
    Generic Library         	                          �         ~�         ~�    �         ��         ��    �         ��         ��    �         �         �    �         ��         ��    �         �         �    �         >�         >�    �         A                             Generic Library         	                         �   	      F         F    �   
      �         �    �         b�         b�    �         �         �    �         V
         V
    �         ��         ��    �                      �       B                            
 LS Library	                �         �    �         �m         �m    �         �N         �N    �          �          �    �         �         �    �   	      2�         2�    �   
      |�         |�    �         �         �    �                      �         R�         R�    �         v         v    �         �5         �5    �         N          N     �         ��         ��    �                �� H��C 4-BITFA2.CKT C:\CIRCUITS\4-BITFA2.CKT 4-BITFA2.CKTA w ���    B w ���   C-in  ���   Sum   ���    C-out ���   ����������������������������  �� �� �� �� �� �� �� �� ��
 �� �� �� �� ��  ���� 
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ���� `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                            ��     ��        ��       ��       ��       ��       ��       ��       ��           ��  	          
     ��                  ��                 ��        ��       ��   
 LS Library	               .P         .P    �         �         �    �         �          �     �         ƚ         ƚ    �         r         r    �                      �         @�         @�    �         �         �    �         jv         jv    �         �o         �o    �         b�         b�    �         �p         �p    �         ��         ��    �         �         �    �         	   
    �� H��C 4-BITFA2.CKT C:\CIRCUITS\4-BITFA2.CKT 4-BITFA2.CKTA out ���    B out ���   C-in  ���   Sum   ���    C-out ���   ����������������������������  �� �� �� �� �� �� �� �� ��
 �� �� �� �� ��  ���� 
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ���� `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                            ��     ��        ��       ��       ��       ��       ��       ��       ��           ��  	          
     ��                  ��                 ��        ��       ��   `
 LS Library               ��         ��    �         ^�         ^�    �         b�         b�    �         {         {    �         n�         n�    �         �         �    �         ΐ         ΐ    �         ~�         ~�    �          .�         .�    �         ރ         ރ    �         �         �    �         ��         ��    �         �v         �v    �         �r         �r    �         Nn         Nn    �         ��         ��    �           ��                                                `
 LS Library              ^�         ^�    �   	      �>         �>    �   
      8�         8�    �         �         �    �         v.         v.    �         ��         ��    �         t�         t�    �         �         �    �         f         f    �   	      �         �    �   
      ��         ��    �         f         f    �                      �         V&         V&    �         $         $    �         �#         �#    �          ��                                                
 LS Library         	                         �        C-in                         `
 LS Library       ,        �7         �7    �         :5         :5    �         �4         �4    �         ><         ><    �         �9         �9    �         �9         �9    �         @         @    �         �?         �?    �         ��         ��    �         T�         T�    �         ��         ��    �         `�         `�    �         V         V    �         *1         *1    �         �0         �0    �         �-         �-    �          !  ��                                                
 LS Library         /        H�         H�    �         ��         ��    �         h�         h�    �         ��         ��    �         V          V     �         ZM         ZM    �         
M         
M    �         >C         >C    �   !     Sum                          	 
 LS Library         /        2�         2�    �   $     C-out                                                                                                               	        
                                                                                                                                         	                                  	   
  	                              "  "   
 #    #   $ % %                                           	 
                                 	 
              &               &                                       	        
   
 &               &                                                     	 
                                                                        (          (                	         	 
             	 
            	 
                              	            	                   ,                ,             ! /                      " ,            # ,            $ /   	                   A      B     C-in     Sum   	  C-out 	                     P xd       �An                                                        