     :
 LS Library       $                          �         �,         �,    �         F,         F,    �         6  ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �         7  ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��      
 LS Library                                  �   	     C-in                         
 LS Library                                  �   
     Y                            
 LS Library                                   �        X                            :
 LS Library       -                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��      
 LS Library         O        �k         �k    �   4      C-out                         
 LS Library         O  
      g         g    �   5     Sum                                                                                                      
         
             
                  	    	      	   
  	                  , ,            $   7              	   
 
                     6     $  $ %  % !  # &  ' &  '    (  ( )  )    *  + *  +   & ,  ,    	 - !  - " . - # . " $ , 2 % 2 / &  3 ' 3 0 (   5 ) 1 4 *    +   8 8   * 
    *     $             $ 	             *          $           $            !                                   	             
         
     	       	     -            -       +    2            *      *    *     +     #           #           #       &          
                	     	                 @            @           E            @            @       !    E          	  H   	         H   	      	   M   	     (  
 ! 8   
        " 8   
    #   # =   
        $ 6          % 6         & ?          ' ?         ( F         ) F         * F        	 + F        	 , ?       $   - 6     !   "   . 6     " #   / @        %   0 @       '   1 E        )   2 ?     $ %   3 #     & '   4 O        )   5 O        (  
 6 ) 
           7 )               0  D   Full Adder       C-out     C-in     Y     X     Sum                      P xd      �An                                                        