     
 LS Library                                   �          A                            
 LS Library                                  �        B                            
 LS Library                                  �        C                            
 LS Library          $                        �        D                            =
 LS Library       $                          �         ��         ��    �        ��      =
 LS Library       $                         �         �T         �T    �        ��      =
 LS Library       $                         �         �3         �3    �      	  ��      =
 LS Library       $ $                        �         ^         ^    �   
     ��      D
 LS Library       0                         �         �         �    �         b�         b�    �         �         �    �              ��      	 D
 LS Library       0                         �         ��         ��    �         ��         ��    �   	      B�         B�    �              ��      
 D
 LS Library       0                         �         ��         ��    �         ^7         ^7    �   
      �"         �"    �              ��       D
 LS Library       0 $                        �         Z�         Z�    �          i         i    �         *g         *g    �              ��       H
 LS Library       0 ,                        �         �j         �j    �         �         �    �         �j         �j    �         �l         �l    �                  ��"       M
 LS Library       8 (                        �         |r         |r    �         lC         lC    �   !   "   #  ��(       M
 LS Library       8                         �   	      &{         &{    �         ��         ��    �   $   %   &  ��(       M
 LS Library       @                         �   
      .�         .�    �         �         �    �   '   (   )  ��(       M
 LS Library       H                         �         ��         ��    �         �         �    �   0   1   2  ��(       
 LS Library         O                         �   3     d                                                                    	                             	              	   
              
               
                	  	       
  
                                                                 < <    6   H    8   K   *  * $  +   + %  & , 	 , ' 
 -   - (   .  . !  /    / "  2 3  ) 4  4 0  5 #  5 1   :   6  @   7    8  9   B C   :  : ;  ;    <   = @ ! =  " 6 ? # < = $ 7 ? % ?  & 	 > ' > A ( A  ) B  * 9 B +  C , 8 D - D  . @ E / E  0 A F 1 F  2 ; G 3 G  4  H 5 H I 6 I  7 F J 8 J  9 
 K : K L ; L  M M                                           %           $             )            $        4    )            $           	 )        &   
 $ %       9    ) %       +    0           0            0           5            0   	         0   	    !    0   	    %    5   	       	  0   
         0   
    (    0   
    )    5   
     
  
  0 %       /    0 &      1    0 '      -     5 &           0 -       3    0 .      6    0 0      8    0 1      ;     5 /          ! 8 )          " 8 +         # = *          $ 8           % 8         	 & =           ' @        	   ( @         
 ) E           * 5         + 5        	 , =      	   - 5     
   
 . 5 )        / 5 +        0 H           1 H          2 M           3 O           4 E         5 =         6 !        "   7 !      $   8 #       ,    9 ,     *    : /          ; /       2   < .      #   = .     ! #     > -     & '   ? !     % $ "   @ .        .   A -     ( ' 0   B ,     ) *    C , %    +    D # '    , -    E . %    . /   F - &    1 0 7   G / -    2 3   H "     4  5   I " .    5 6   J - 0    7 8   K   %    9  :   L   1    : ;       !  5   7-SEGMENT DISPLAY (d)        A      B     C     D     d                      P xd       �An                                                        