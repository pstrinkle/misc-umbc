     
 LS Library	  	     ! 	        ��         ��    �         �]         �]    �         lm         lm    �         m         m    �         
F         
F    �         ��         ��    �         b�         b�    �         ��         ��    �         �         �    �   	      �*         �*    �   
      &�         &�    �         ��         ��    �         F�         F�    �         
         
    �                               	  
        �� |��C 4-BITFA.CKT C:\4-BITFA.CKT 4-BITFA.CKTa1  �V�    b1  �V�   a2  �V�   b2  �V�   a3  �V�   b3  �V�   a4  �V�  	 b4  �V�  
 C-in1 �V�   S1 n1 �V�    S2 n1 �V�   S3 n1 �V�   S4 n1 �V�   C-out4 V�   ���������������������������� �� �� �� ��
 ��	 �� �� �� �� �� �� �� �� ��    
 LS Library                6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                 �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �         ޗ         ޗ    �         t�         t�    �          ��         ��    �         �>         �>    �              	  �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �   	      ޗ         ޗ    �   
      t�         t�    �         ��         ��    �         �>         �>    �   
             �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library        "       6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ����������������������������                    ��        ��                   ��        ��       ��       ��        ��   	     ��  
     ��                 ��       ��       ��        ��       ��  �� 
 LS Library         . 
 	                       �         S1                           �� 
 LS Library         .  
                       �         S2                            
 LS Library         .                         �        S3                            
 LS Library         .                         �        S4                            
 LS Library         /                         �        S5                            
 LS Library         /                          �   "     S6                           	 
 LS Library         / "                        �   #     S7                           
 
 LS Library         / $                        �   $     S8                            
 LS Library         / &                        �   %   	  C-out                         
 LS Library          
                         �   &  
   a1                           
 LS Library                                  �   '     b1                           
 LS Library                                  �   (     a2                           
 LS Library                                  �   )     b2                           
 LS Library                                  �   @     a3                           
 LS Library                                  �   +     b3                           
 LS Library                                  �   ,     a4                           
 LS Library                                  �   -     b4                           
 LS Library          ,                        �   V     b8                           
 LS Library          *                        �   W     a8                           
 LS Library          (                        �   X     b7                           
 LS Library          &                        �   Y     a7                           
 LS Library          $                        �   Z     b6                           
 LS Library          "                        �   [     a6                           
 LS Library                                   �   \     b5                           
 LS Library	  	     "        ��         ��    �         �]         �]    �         lm         lm    �         m         m    �         
F         
F    �         ��         ��    �         b�         b�    �         ��         ��    �         �         �    �         �*         �*    �         &�         &�    �         ��         ��    �         F�         F�    �         
         
    �   5   4   3   2   1   0   /   .                �� |��C 4-BITFA.CKT C:\4-BITFA.CKT 4-BITFA.CKTa1  O�    b1  O�   a2  O�   b2  O�   a3  O�   b3  O�   a4  O�  	 b4  O�  
 C-in1 O�   S1 n1 O�    S2 n1 O�   S3 n1 O�   S4 n1 O�   C-out4 �   ���������������������������� �� �� �� ��
 ��	 �� �� �� �� �� �� �� �� ��    
 LS Library                6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                 �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �         ޗ         ޗ    �         t�         t�    �          ��         ��    �         �>         �>    �              	  �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �   	      ޗ         ޗ    �   
      t�         t�    �         ��         ��    �         �>         �>    �   
             �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library        "       6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ����������������������������                    ��        ��                   ��        ��       ��       ��        ��   	     ��  
     ��                 ��       ��       ��        ��       ��   
 LS Library                                  �   6     C-in                         
 LS Library                                  �        a5                                                                                                                        	           
                                                                                                                                        	         
             J H   6 7  7 8  8   & :  : 9  >   <   ( ;  < ; 	 '  
 ) =  > =  9    * ?  @ ?  *   + A  B A  B   , C  D C  D   - E  F E  F   s k  t l  u m �� w o  x p  q y   
 h ! f  ��# V k $ W l % v n & X m ' Y n (  q ) i  * s . + t / , u 0 - v 1 . w 2 / x 3 0 Z o 1 y 5 2 j i 3 j r 4  r 5 	  6 g f 7  g 8 h   9  e : e d ; d  <   =  b > b " ?  c @ c a A a # B  ` C ` _ D _ $ E  ^ F ^ ] G ] % H [ p I \ 4 z c   !              !        	    !            !            !            !            !            !            !           	 )         5  	 
 )           
  )        7    )        9    )        4   ��������������         (    * #      E    * "      B    * !      ?    *        =    *        <    "       )    .        5  	  /        <    .        ;    .        !     .        8  
 ��" / !       >   # / #  	     A   $ / %  
     D   % / '       G   &             '         	   (            )         
   *          +            ,            -            . " '      *   / " &      +   0 " %      ,   1 " $      -   2 " #      .   3 " "      /   4 " !      I   5 "         1   6  	           7  	         8          9           :           ;          <          =      
    >          ?          @            A          B          C          D          E           F           ������������������������������V  -       #   W  +       $   X  )       &   Y  '       '   Z  %       0   [  #       H   \  !       I   ] , '    F G   ^ , #    E F   _ - %    C D   ` - "    B C   a . #    @ A   b /      = >   c . !    ? @   d ,     : ;   e ,     9 :   f -     6 !   g -     7 6   h .     8    
 i       2 )   j       3 2   k ! -     #   l   +     $   m  )     &   n  '    % '   o  %     0   p  #     H   q       (   r )     4 3   s ! '    *    t   &    +    u  %    ,    v  $    - %   w  #    .    x  "    /    y       1              S1  ��   S2     S3     S4     S5     S6   	  S7 	  
  S8 
 	   C-out  
   a1     b1     a2     b2     a3     b3     a4     b4  ��   b8     a8     b7     a7     b6     a6     b5     C-in     a5                              	 	  
 
                                                   P xd       �An                                                        