      Generic Library                                   �                      �         0�         0�    �         \�         \�    �         A                             Generic Library         
                         �         `�         `�    �         ��         ��    �         T�         T�    �       B                            
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  љo    Y in  љo   X in  љo   C-out љo    Sum t љo   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  љo    Y in  љo   X in  љo   C-out љo    Sum t љo   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  љo    Y in  љo   X in  љo   C-out љo    Sum t љo   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  љo    Y in  љo   X in  љo   C-out љo    Sum t љo   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library         /  
      ��         ��    �         B�         B�    �         ��         ��    �         ��         ��    �        Sum                           
 LS Library         /        ��         ��    �        C-out                         `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                             
 LS Library                                  �   5     C-in                                                                                                           	          
                                                               5 5    %  %     $  $ &  & !  '   ' "   (  ) ( 	 ) # 
  *  + *  +    ,  . ,  . -  
 /  -   0 /  0 1  1    2  3 2  3 4  4   5 6  6 7  7    8   9  :   : 9     ! 8 ; " ; < # < 	 $  = % = > & >  '  ? ( ? @ ) @ A * A B + B  ,  C - C D . D  /  E 0 F  1 G F 2  G 3 E H 4 H  I I    	                           	                           
            	            ( 
         	  ( 	         
             	          .   	         #   
 (            (                                0            &    (            (             "             !      4             +    ( !       
    (            /       
       
     /             	              
                 $           '       	            	    ,       	    2       	    /     ,   
       
 ! ,   
       " ,   
       # ,   
    	   $ +         % , 	        
 & +         ' (         ( )          ) )      	   * * !    
    + *         , (         -  "        .          / (         0          1          2 (        	 3         	 4         	 5            6          7          8  
     !   9          :  
        ;      ! "   <       " #   =      $ %   >      % &   ?      ' (   @      ( )   A      ) *   B       * +   C      , -   D      - .   E      / 3   F      1 0   G      2 1   H  !    3 4              A      B     Sum     C-out     C-in                      P xd       �An                                                        