     
 LS Library                                   �          A                            
 LS Library                                  �        B                            
 LS Library                                  �        C                            
 LS Library                                  �        D                            s
 LS Library         9                         �         &{         &{    �         �~         �~    �         lC         lC    �         |r         |r    �   	      �,         �,    �   
      �l         �l    �                  	   
   ��  
 LS Library       '         �}         �}    �         �j         �j    �         �         �    �         �j         �j    �         �          �     �                 �� ��C
 7SEG-A.CKT C:\7SEG-A.CKT
 7SEG-A.CKTA � �2G    B � �2G   C � �2G   D � �2G   a � �2G    ����������  �� �� �� �� ��  �������� =
 LS Library                                  �         B�         B�    �        ��      =
 LS Library                                 �         B�         B�    �        ��      =
 LS Library                                  �         �T         �T    �      	  ��      =
 LS Library         (                        �         ��         ��    �   
     ��      A
 LS Library       ,                         �         Ɛ         Ɛ    �         r�         r�    �           ��      	 D
 LS Library       ,                         �         �         �    �         j�         j�    �   	      �3         �3    �              ��      
 D
 LS Library       ,                          �         �/         �/    �         "�         "�    �   
      Z�         Z�    �              ��       D
 LS Library       ,                          �         *g         *g    �         �          �     �         �j         �j    �              ��       M
 LS Library       4                         �         �l         �l    �         �j         �j    �   -   .   /  ��(       M
 LS Library       4  	                       �   
      �l         �l    �         �,         �,    �   0   1   2  ��(       M
 LS Library       =                         �         |r         |r    �         lC         lC    �   3   4   5  ��(      ��     ��             ��      	     ��           ��      	             	             
             
         
            	  	        
  
                                          ��    
 LS Library       '        z�         z�    �         @z         @z    �         z@         z@    �          ��         ��    �         08         08    �                 �� �C
 7SEG-B.CKT C:\7SEG-B.CKT
 7SEG-B.CKTD � �2G    C � �2G   B � �2G   A � �2G   b � �2G    ����������  �� �� �� �� ��  ���������� =
 LS Library        (                         �         b�         b�    �        ��      =
 LS Library                                 �         b�         b�    �        ��      =
 LS Library                                �         ��         ��    �   	   
  ��      =
 LS Library                                �         ^         ^    �        ��     	 A
 LS Library       '                         �         r�         r�    �         ��         ��    �           ��      
 D
 LS Library       '                         �         j�         j�    �         �3         �3    �   	      �1         �1    �              ��       D
 LS Library       '                          �         "�         "�    �          Z�         Z�    �   
      i         i    �              ��       D
 LS Library       '                         �         �          �     �         �j         �j    �         �         �    �              ��       M
 LS Library       0  	                       �   
      ��         ��    �         �j         �j    �           ��(       M
 LS Library       0                         �         �,         �,    �         z.         z.    �          !  ��(       M
 LS Library       8                         �         lC         lC    �         �~         �~    �   "   #   $  ��(      ��     ��            ��           ��        ��                
         
            	            	    
          	       	  
        
                                            ��    
 LS Library       '        p�         p�    �         ܭ         ܭ    �         ��         ��    �          ��         ��    �         B�         B�    �                 �� ��C
 7SEG-C.CKT C:\7SEG-C.CKT
 7SEG-C.CKTD � �2G    C � �2G   B � �2G   A � �2G   c � �2G    ����������  �� �� �� �� ��  �������� =
 LS Library        $                         �         �,         �,    �        ��      =
 LS Library                                �         �j         �j    �        ��     �� =
 LS Library                                �         �j         �j    �   
     ��      =
 LS Library                                �         *g         *g    �        ��     	 A
 LS Library       (                         �         Z�         Z�    �         "�         "�    �           ��      
 A
 LS Library       (                         �          �1         �1    �   	      �3         �3    �           ��       D
 LS Library       (                         �         �         �    �         ��         ��    �   
      r�         r�    �              ��       D
 LS Library       ( $                        �         ^         ^    �         ��         ��    �         ��         ��    �              ��       M
 LS Library       0   
                       �         b�         b�    �         �         �    �           ��(       M
 LS Library       0                         �   	      �         �    �         B�         B�    �          !  ��(       M
 LS Library       8                         �         ��         ��    �         B�         B�    �   "   #   $  ��(      ��     ��       
     ��        ��      	     ��                                                  	    
      	        	  
       
                                            ��    
 LS Library       '         0M         0M    �         <         <    �         ��         ��    �         ^�         ^�    �         "{         "{    �                 �� ��C
 7SEG-D.CKT C:\7SEG-D.CKT
 7SEG-D.CKTA � �2G    B � �2G   C � �2G   D � �2G   d � �2G    ����������  �� �� �� �� ��  �������� =
 LS Library       $                          �         ��         ��    �        ��      =
 LS Library       $                         �         �T         �T    �        ��      =
 LS Library       $                         �         �3         �3    �      	  ��      =
 LS Library       $ $                        �         ^         ^    �   
     ��      D
 LS Library       0                         �         �         �    �         b�         b�    �         �         �    �              ��      	 D
 LS Library       0                         �         ��         ��    �         ��         ��    �   	      B�         B�    �              ��      
 D
 LS Library       0                         �         ��         ��    �         ^7         ^7    �   
      �"         �"    �              ��       D
 LS Library       0 $                        �         Z�         Z�    �          i         i    �         *g         *g    �              ��       H
 LS Library       0 ,                        �         �j         �j    �         �         �    �         �j         �j    �         �l         �l    �                  ��"       M
 LS Library       8 (                        �         |r         |r    �         lC         lC    �   !   "   #  ��(       M
 LS Library       8                         �   	      &{         &{    �         ��         ��    �   $   %   &  ��(       M
 LS Library       @                         �   
      .�         .�    �         �         �    �   '   (   )  ��(       M
 LS Library       H                         �         ��         ��    �         �         �    �   0   1   2  ��(      ��     ��            ��           ��      	        ��                   	              	   
              
               
                	  	       
  
                                                             ��   	 
 LS Library       '          Z�         Z�    �         :X         :X    �         �m         �m    �         *b         *b    �         2^         2^    �          !   "   #  �� ��C
 7SEG-E.CKT C:\7SEG-E.CKT
 7SEG-E.CKTA � �2G    B � �2G   C � �2G   D � �2G   e � �2G    ����������  �� �� �� ��
 ��  �������� =
 LS Library         $                        �         ��         ��    �        ��      =
 LS Library                                 �         B�         B�    �        ��      =
 LS Library                                 �         b�         b�    �      	  ��      =
 LS Library                                  �         b�         b�    �   
     ��      D
 LS Library       ,                         �         ��         ��    �         ��         ��    �         ^         ^    �              ��      	 D
 LS Library       ,                         �         r�         r�    �         ��         ��    �   	      �         �    �              ��      
 M
 LS Library       9                         �   	      �3         �3    �   
      �1         �1    �           ��(      ��     ��         ��           ��        ��               	         	         	                    
    	  	    
   
  
    ��   
 
 LS Library       ' &        d�         d�    �         @�         @�    �         ��         ��    �         Y         Y    �   	      �a         �a    �   $   %   &   '   (  �� �	�C
 7SEG-F.CKT C:\7SEG-F.CKT
 7SEG-F.CKTA � �2G    B � �2G   C � �2G   D � �2G   f � �2G    ����������  �� �� �� �� ��  �������� =
 LS Library       $ $                        �         ��         ��    �        ��      =
 LS Library       $                         �         Ɛ         Ɛ    �        ��      =
 LS Library       $                         �         ��         ��    �      	  ��      =
 LS Library       $                          �         �T         �T    �   
     ��      D
 LS Library       0                         �         �         �    �         b�         b�    �         �         �    �              ��      	 D
 LS Library       0                         �         ��         ��    �         ��         ��    �   	      B�         B�    �              ��      
 D
 LS Library       0                         �         ��         ��    �         ^7         ^7    �   
      �"         �"    �              ��       D
 LS Library       0 $                        �         Z�         Z�    �          i         i    �         *g         *g    �              ��       M
 LS Library       8                         �   	      �j         �j    �         �         �    �   -   .   /  ��(       M
 LS Library       8   
                       �         �l         �l    �         �,         �,    �   0   1   2  ��(       M
 LS Library       @                         �         lC         lC    �         �~         �~    �   3   4   5  ��(      ��     ��            ��         
     ��        ��            	   
            	                          	    
              	  	       
  
                                          ��    
 LS Library       ' ,                     �         B�         B�    �         ��         ��    �         J�         J�    �   
      p6         p6    �   )   *   +   ,   -  �� �
�C
 7SEG-G.CKT C:\7SEG-G.CKT
 7SEG-G.CKTA � �2G    B � �2G   C � �2G   D � �2G   g � �2G    ����������  �� �� �� �� ��  �������� =
 LS Library       $ $                        �         ��         ��    �        ��      =
 LS Library       $                         �         �~         �~    �        ��      =
 LS Library       $                         �         |r         |r    �      	  ��      =
 LS Library       $                          �         �l         �l    �   
     ��      D
 LS Library       0                         �         �         �    �         �j         �j    �         �          �     �              ��      	 D
 LS Library       0                         �         i         i    �         Z�         Z�    �   	      "�         "�    �              ��      
 D
 LS Library       0                         �         ^7         ^7    �         ��         ��    �   
      B9         B9    �              ��       D
 LS Library       0 $                        �         ��         ��    �          ��         ��    �         B�         B�    �              ��       M
 LS Library       8                          �         b�         b�    �         �         �    �   -   .   /  ��(       M
 LS Library       8  
                       �   	      ^         ^    �         Ɛ         Ɛ    �   0   1   2  ��(       M
 LS Library       @                         �         XU         XU    �          �          �    �   3   4   5  ��(      ��     ��            ��        ��      	   
     ��            
                     	                
    	                  	  	       
  
                                          ��                           
        	                      
      	                     
      	                       
      	                                             	    	     
    
         S S    .  . /  /   0   0    1  2 1   3  2  	 4 3 
 4   # 5  6 5  6   ( 7  8 7  8 	  - 9  : 9  : 
  ;    ; B   <  = <  = D   >  ? >  ? F   @  A @  A H   B   B C ! C  "  D # D E $ E  %  F & F G ' G  (  H ) H I * I  + C J , J  - E K . K  / G L 0 L  1 I M 2 M  3 J N 4 N  5 K O 6 O  7 L P 8 P  9 M Q : Q  ; N R < R  = O S > S   ? P T @ T ! A Q U B U " C R V D V $ E S W F W % G T X H X & I U Y J Y ' K V Z L Z ) M W [ N [ * O X \ P \ + Q Y ] R ] , c ^                                                     9            9           9           9       
    9          	 9         	 
 9         
  ' 
            '       "    '       %    '       (    / 
            '        2    /            '       !     '       $    '       '    '        *    '       0    '       .    '       ,     /            '        4     '       6    '       8    '       :    /            ' "  	     <      ' #  	    >   ! ' $  	    @   " ' %  	    B   # / "  	        $ ' (  
     D    % ' )  
    F   & ' *  
    H   ' ' +  
    J   ( / (  
       	 ) ' .       L    * ' /      N   + ' 0      P   , ' 1      R   - / .         
 . 8 
         / 8         0 /         1 0         2 0         3 1      	   4 1     	 
   5 2 "        6 2         7 3 (       	 8 3        	 9 4 .       
 : 4        
 ;  
         <          =          >          ?          @          A          B & 
           C &     !   +    D %     "  #   E %     $ # -   F $     %  &   G $     ' & /   H #     (  )   I #     * ) 1   J &     , + 3    K %     . - 5   L $     0 / 7   M #     2 1 9   N &     4 3 ;    O %     6 5 =   P $     8 7 ?   Q #     : 9 A   R & "    ; C <    S % #    = E >   T $ $    ? G @   U # %    A I B   V & (    D C K    W % )    F E M   X $ *    H G O   Y # +    J I Q   Z & .    K L    [ % /    M N   \ $ 0    O P   ] # 1    Q R   ����������    !  5   7-SEGMENT DISPLAY        A      B     C     D                   P xd       �An                                                        