     
 LS Library 	      $         &          &     �         ��         ��    �         J�         J�    �         ��         ��    �         ��         ��    �         V�         V�    �         �         �    �         N�         N�    �         �u         �u    �   	      l         l    �   
      �         �    �         �<         �<    �         ��         ��    �          V          V    �         r�         r�    �         �         �    �         �         �    �         ��         ��    �         ��         ��    �         ��         ��    �         �"         �"    �         Đ         Đ    �         �P         �P    �         r�         r�    �         ҥ         ҥ    �         &�         &�    �                 �� ��C 8-BITFA2.CKT C:\CIRCUITS\8-BITFA2.CKT 8-BITFA2.CKTA � �V�    B � �V�   C-in  �V�   Sum   �V�    C-out �V�   ����������������������������������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��
  ���� 
 LS Library	                �         �    �         �m         �m    �         �N         �N    �          �          �    �         �         �    �   	      2�         2�    �   
      |�         |�    �         �         �    �                      �         R�         R�    �         v         v    �         �5         �5    �         N          N     �         ��         ��    �                �� H��C 4-BITFA2.CKT C:\CIRCUITS\4-BITFA2.CKT 4-BITFA2.CKTA � �V�    B � �V�   C-in  �V�   Sum   �V�    C-out �V�   ����������������������������  �� �� �� �� �� �� �� �� ��
 �� �� �� �� ��  ���� 
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ���� `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                            ��     ��        ��       ��       ��       ��       ��       ��       ��           ��  	          
     ��                  ��                 ��        ��       ��   
 LS Library	               .P         .P    �         �         �    �         �          �     �         ƚ         ƚ    �         r         r    �                      �         @�         @�    �         �         �    �         jv         jv    �         �o         �o    �         b�         b�    �         �p         �p    �         ��         ��    �         �         �    �         	   
    �� H��C 4-BITFA2.CKT C:\CIRCUITS\4-BITFA2.CKT 4-BITFA2.CKTA out �V�    B out �V�   C-in  �V�   Sum   �V�    C-out �V�   ����������������������������  �� �� �� �� �� �� �� �� ��
 �� �� �� �� ��  ���� 
 LS Library                2�         2�    �         ��         ��    �          �.         �.    �   	      b*         b*    �   
      �
         �
    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library          	                     �         ��         ��    �         H;         H;    �         �         �    �         t         t    �         	   
    �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                Z�         Z�    �         @2         @2    �         v�         v�    �         �         �    �         �         �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                �         �    �         ��         ��    �         ^�         ^�    �         ��         ��    �          �          �    �                �� ���C FA.CKT C:\CIRCUITS\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ���� `
 LS Library       	        2�         2�    �         .         .    �         b]         b]    �         �-         �-    �          �?         �?    �         �?         �?    �         �         �    �         �         �    �               ��
                                            	 `
 LS Library              �         �    �         >         >    �         �         �    �         �         �    �         C         C    �         �B         �B    �         VQ         VQ    �         Q         Q    �              ��
                                            
 `
 LS Library       ,  
      �V         �V    �         �V         �V    �         �^         �^    �         �^         �^    �   
      �E         �E    �         NE         NE    �         �g         �g    �         Dg         Dg    �       !   "   #     ��                                            ��     ��        ��       ��       ��       ��       ��       ��       ��           ��  	          
     ��                  ��                 ��        ��       ��   `
 LS Library               ��         ��    �         ^�         ^�    �         b�         b�    �         {         {    �         n�         n�    �         �         �    �         ΐ         ΐ    �         ~�         ~�    �          .�         .�    �         ރ         ރ    �         �         �    �         ��         ��    �         �v         �v    �         �r         �r    �         Nn         Nn    �         ��         ��    �           ��                                                `
 LS Library              ^�         ^�    �   	      �>         �>    �   
      8�         8�    �         �         �    �         v.         v.    �         ��         ��    �         t�         t�    �         �         �    �         f         f    �   	      �         �    �   
      ��         ��    �         f         f    �                      �         V&         V&    �         $         $    �         �#         �#    �          ��                                               �� `
 LS Library       ,        �7         �7    �         :5         :5    �         �4         �4    �         ><         ><    �         �9         �9    �         �9         �9    �         @         @    �         �?         �?    �         ��         ��    �         T�         T�    �         ��         ��    �         `�         `�    �         V         V    �         *1         *1    �         �0         �0    �         �-         �-    �          !  ��                                               ����     ��         ��       ��       ��       ��        ��       ��       ��       ��     	  �� 	    
  �� 
      ��       ��       ��       ��       ��          ��        ��        ��       ��       ��                ��       ��       ��       ��       ��  ������ 
 LS Library                                   �         �         �    �         ��         ��    �         B�         B�    �         ��         ��    �         F�         F�    �         ��         ��    �         ��         ��    �   	    A                            
 LS Library                                  �   
     C-in                         
 LS Library                                  �         "         "    �         �9         �9    �         �=         �=    �         @A         @A    �          E          E    �          �         �    �   !      F         F    �   l    B                            
 LS Library         0        ��         ��    �         �         �    �         n�         n�    �         ��         ��    �         ʖ         ʖ    �         ��         ��    �         z�         z�    �         j�         j�    �        Sum                           
 LS Library         0        چ         چ    �        C-out                        �������������������������������� 
 LS Library	               �         �    �         D�         D�    �         vc         vc    �         �b         �b    �         6b         6b    �         �a         �a    �          �`         �`    �   !      V`         V`    �         zB         zB    �         >;         >;    �   	      �:         �:    �   
      &C         &C    �         F@         F@    �         �?         �?    �         ?         ?    �         �_         �_    �         _         _    �      k   j  �� 6��C 8-BITXOR.CKT C:\CIRCUITS\8-BITXOR.CKT 8-BITXOR.CKTB � �V�    C-in  �V�   XOR'd �V�    ����������������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� 
 ���� ]
 LS Library                                  �         t�         t�    �   	      $�         $�    �           ��3        ]
 LS Library                                 �         ��         ��    �   
      ��         ��    �           ��3        ]
 LS Library                                 �         D�         D�    �         �         �    �      	   
  ��3        ]
 LS Library         %                        �         �y         �y    �         By         By    �           ��3        ]
 LS Library         +                        �         �k         �k    �         �k         �k    �           ��3        ]
 LS Library         0                        �         .^         .^    �         �]         �]    �           ��3        ]
 LS Library         6                        �         |P         |P    �         ,P         ,P    �           ��3       	 ]
 LS Library         ;                        �         �B         �B    �         zB         zB    �           ��3       
 `
 LS Library               8�         8�    �         �         �    �         �I         �I    �         �I         �I    �         >I         >I    �         �H         �H    �         �H         �H    �         NH         NH    �          �G         �G    �         �G         �G    �         ^G         ^G    �         G         G    �         �F         �F    �         nF         nF    �         F         F    �         �E         �E    �                  !      ��                                                                                 `
 LS Library       0  	      �D         �D    �   
      �B         �B    �         ~B         ~B    �         .B         .B    �         �A         �A    �         �A         �A    �         >A         >A    �         �@         �@    �   	      �@         �@    �   
      N@         N@    �         �?         �?    �         �?         �?    �         ^?         ^?    �         ?         ?    �         �>         �>    �         n>         n>    �   9   :   ;   <   =   >   ?   @   A  ��                                                                                ��     ��         ��        ��        ��        ��        ��        ��        ��  	     	 ��                       	   	      ��   
      ��        ��        ��        ��        ��        ��    	    ��  " "                                                                                      	     	    
     
                                                                                                                                                                                                             !        N  ������            ��   ����������������������������������������������������������������������������������������������������������������������D f  E 	 f F    G g  H g h I  i J i k K j h L l  M 
 i m    $         F            $        G   	 
       $            ,                    ,           ��������	         E           
  	       M            L          !       F D            0                   0           �� ,           	     I             ����������������������������������������������������������������������������������������������������������������������������������������������������������������������f      E D           g "     H G   	 
      h "     K H   	 
      i  	    J M I   j         K   	 
      k        J   l         L          !       ����   A     C-in     B     Sum     C-out                    P xd       �An                                                        