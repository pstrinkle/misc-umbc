     
 LS Library                6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                 �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �         ޗ         ޗ    �         t�         t�    �          ��         ��    �         �>         �>    �              	  �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �   	      ޗ         ޗ    �   
      t�         t�    �         ��         ��    �         �>         �>    �   
             �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library        "       6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library                                  �         a1                           
 LS Library                                  �        b1                           
 LS Library                                  �        a2                           
 LS Library                                  �        b2                           
 LS Library           
                       �        a3                          	 
 LS Library           	                       �        b3                          
 
 LS Library          "                        �        a4                           
 LS Library          $                        �        b4                           
 LS Library         (                         �        S1                            
 LS Library         (                         �      	  S2                            
 LS Library         (                         �      
  S3                            
 LS Library         ( #                        �        S4                            
 LS Library         ( &                        �         C-out4                        
 LS Library          
                        �   - 	    C-in1                                                                                                                   	     	    
                                          
                       ) )   # "   #  ! "  ! $  $     %  % &  ' &  ' ( 	 ( 
 
  )  ) *  + *  + ,  ,   - .  . /  /    0  0 1  1          2  2 3  3    4  4 5  5      7 6   7     ! 6  " 	  #   $   %   &  8 ' 8 9 ( 9   : :                                         $             $        #                                      $            	 $       "   
         	             	           
  $        
    $       $     &            %            $      !    $ %       &    $ $      %                                                              
     	       	   #  
          %            (        "    (        #    (        $    ( $       %     ( '       (   !           " %           # %           $           % %         & %         '          (       	   ) %     
    * % !        +  !        ,  &        -            .          /          0          1          2          3          4         
 5         
 6  $     !   7  #        8 & %    & '   9 & '    ' (         0   4-bit Adder       a1     b1     a2     b2     a3   	  b3 	  
  a4 
    b4     S1  	   S2  
   S3     S4     C-out4     C-in1                                 	 	  
 
            P xd       �An                                                        