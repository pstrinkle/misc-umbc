   �� 
 LS Library          (                         �        D                            
 LS Library                                   �        C                            
 LS Library                                  �        B                            
 LS Library                                  �        A                            =
 LS Library        (                         �         b�         b�    �        ��      =
 LS Library                                 �         b�         b�    �        ��      =
 LS Library                                �         ��         ��    �   	   
  ��      =
 LS Library                                �         ^         ^    �        ��     	 A
 LS Library       '                         �         r�         r�    �         ��         ��    �           ��      
 D
 LS Library       '                         �         j�         j�    �         �3         �3    �   	      �1         �1    �              ��       D
 LS Library       '                          �         "�         "�    �          Z�         Z�    �   
      i         i    �              ��       D
 LS Library       '                         �         �          �     �         �j         �j    �         �         �    �              ��       M
 LS Library       0  	                       �   
      ��         ��    �         �j         �j    �           ��(       M
 LS Library       0                         �         �,         �,    �         z.         z.    �          !  ��(       M
 LS Library       8                         �         lC         lC    �         �~         �~    �   "   #   $  ��(       
 LS Library         ?        ��         ��    �   A     b                                                                                       
         
            	            	    
          	       	  
        
                                                2 2   1 2  '   + (   (  ) ,   )  . 4  % /  0 - 	 * 0 
  *  & 1  +   ,   -   .   /   0   1    *  
 2   3   4      	   )   (  '   &   / 3  %    5   5 6 ! 6  "  7 # 8 7 $ 8   % ! 9 & 9 : ' : " (  ; ) ; < * <  +  = , > = - >  .  ? / @ ? 0 @ # 1 $ A B A ��  )             !                                    )            ! )            !           ! !          	            
 !                         !            '   	     
    '   	        ,   	     "    '   
         '   
        '   
        ,   
     (  	  ' !           ' "          ' #           , "       +  
  ' 	           ' 
          '           , 
           0        *  	  0       -  
  5        .    0        !     0       $   ! 5        %   " 8        '   # 8       0   $ =        1   % $         & % 
        '  	        (  )          )  !         * &     
  	   +  #         ,  "        - & !        . #         / $          0 &      	    1 %           2 %          3 $ !        4 # )        5 . 
         6 .       !   7 .     " #   8 .     # $   9 7     % &   : 7     & '   ; /     ( )  	 < /     ) *  	 = / "    + ,  
 > /     , -  
 ? 7     . /   @ 7     / 0   A ?        1         1   7-SEGMENT DISPLAY (b)   ��   D     C     B     A     b                    P xd       �An                                                        