      Generic Library         	                          �         �8         �8    �         f8         f8    �         8         8    �         �7         �7    �         v7         v7    �         &7         &7    �         �6         �6    �         B                             Generic Library                                  �        C-in                         ]
 LS Library                                  �         t�         t�    �   	      $�         $�    �           ��3        ]
 LS Library                                 �         ��         ��    �   
      ��         ��    �           ��3        ]
 LS Library                                 �         D�         D�    �         �         �    �      	   
  ��3        ]
 LS Library         %                        �         �y         �y    �         By         By    �           ��3        ]
 LS Library         +                        �         �k         �k    �         �k         �k    �           ��3        ]
 LS Library         0                        �         .^         .^    �         �]         �]    �           ��3        ]
 LS Library         6                        �         |P         |P    �         ,P         ,P    �           ��3       	 ]
 LS Library         ;                        �         �B         �B    �         zB         zB    �           ��3       
 `
 LS Library               �?         �?    �         ^3         ^3    �         �         �    �         �         �    �         H         H    �         �         �    �         �         �    �         X         X    �                       �         �         �    �         h         h    �                      �         �         �    �         x         x    �         (         (    �         �         �    �                  !      ��                                                                                 `
 LS Library       0  	      �         �    �   
      l         l    �                      �         �         �    �         |         |    �         ,         ,    �         �         �    �         �         �    �   	      <         <    �   
      �         �    �         �         �    �         L         L    �         �         �    �         �         �    �         \         \    �                      �   9   :   ;   <   =   >   ?   @   A  ��                                                                                 
 LS Library         3  	      v'         v'    �   
      �%         �%    �         B%         B%    �         �$         �$    �         �$         �$    �         R$         R$    �         $         $    �         �#         �#    �   A     XOR'd                                                                                                        	     	                          	   	          
                                                        	       > =       "  " #  #    $  $ %  %    &  & ' 	 '  
  (  ( )  )    *  * +  +     ,  , -  -    /  0   1 0  ! 1  / .  .   . 2  2   2 3  3 	  3 4  4   4 5   5  ! 5 6 " 6  # 6 7 $ 7  % 7 8 & 8  '  9 (  B ) C B * C : + 
 D , E D - E ; .  F / G F 0 G < 1  H 2 I H 3 I = 4  K 5 J K 6 J > 7  L 8 M L 9 M ? :  N ; O N ��= O @ Q P           
                                                        %        '  	                           %        (  
               	   "         
 % !       +      &       	      (          % '       .      ,             .           % -       1      1             3      "    % 2       4      7             9      $    % 8       7      <  	           >  	    &    % =  	     :       
           
           
              
           
    
       
            
       !    
       "          #          $          %           &          '  &     	   (      
    )  ,        *          +  1        ,          -  7        .           /          0  <        1          2           3  "         4  (         5  .       !   6  3    " ! #   7  9    $ # %   8  >    % &   9 0        '  	 : 0       *  
 ; 0       -   < 0       0   = 0       3   > 0       6   ? 0       9   @ 0       =   A 3              	 
       B &     ( )  
 C &     ) *  
 D ' !    + ,   E '     , -   F ( '    . /   G (     / 0   H ) -    1 2   I )     2 3   J *     5 6   K * 2    4 5   L + 8    7 8   M +     8 9   N , =    : ;   O ,     ; =   ��           B      C-in     XOR'd                P xd       �An                                                        