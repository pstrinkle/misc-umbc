     u            u Generic Library       #                          �         ��         ��    �         N�         N�    �          ��         ��    �         ��         ��    �         ^�         ^�    �                  ��      �AN        �@N          Meg         �<N1 u           u Generic Library       #                          �         ֪         ֪    �         ��         ��    �          6�         6�    �         �         �    �         ��         ��    �   H  
   	         ��      �AN        �@N          Meg         �<N1  Generic Library                                  �         C                             Generic Library          +                        �   - 
   Clock                         zDN        �CN       Clock  Generic Library                                   �        PE                           Generic Library         8        ��         ��    �        A                              Generic Library         8        ��         ��    �        B                             D Generic Library                                �   	      ��         ��    �         d�         d�    �   
      �         �    �              ��0       D Generic Library                                �         ��         ��    �         p�         p�    �          �          �    �             !  ��0      	 M Generic Library         
                       �         ��         ��    �         ��         ��    �   "   #   $  ��;      
 D Generic Library                                �         ��         ��    �         R�         R�    �         v�         v�    �   )   *   +   ,  ��0       A Generic Library        !                        �         Rw         Rw    �         �v         �v    �      .   /  ��-       A Generic Library        '                        �         �i         �i    �         Vi         Vi    �   0   1   2  ��-       M Generic Library        $                        �         z�         z�    �         f�         f�    �   3   4   5  ��;       M Generic Library                                �         �S         �S    �         �S         �S    �   6   7   8  ��;       = Generic Library       	                         �   	      j%         j%    �   @   A  ��)      = Generic Library       	                         �         j�         j�    �   >   =  ��)      = Generic Library       	 #                        �         b�         b�    �   R   T  ��)                                    	                        
                                                   
                                 
   	         
      	                   	     
                                             O O   , 9  -               % >  K %    	   
           	      &   E   [  B   ' (    (  D B     9 :  : 6  / 3  4 2  < 7  < 5  ; 8  ; 
  & '   D & ! ! G " ? G # ? # $ $  %  C & H  ' C  ( J  ) J " *  E + F E , K X -   . L I / L % 0  I 1 A  2 =  3 @  4 M  5 M N 6 N   7 B O 8 O  9 O P : P 0 ; N Z < Q R = T . >  S ? S U @ V U A W V B W 1 C F X D X Y E Y ) F Q Z G Z * H  [ I [ \ J ] \ K ] ^ L _ ^ M _ ` N ` + a a   )            )         H    &        -     #            #        $    &              )       >    )            &           	 #          
 #           	     3 ' 4     	       %     "       8                 " ,         "          "           & $          4 $          &      - &     4      	      4     
 	     &       
     8            8        *                       1  	         0            (  
                     2            6   !         !   "    	     )  
 #    	    #   $    	     $   %       /    &  
          ' * 
        ( *         )    
     E   *    
    G   +    
    N   ,    
         -  ,          .  $      =   /  #          0  (       :   1  *      B   2  )          3  %          4  '         5  &          6            7            8 !           9           :          ; !         <           =         2   > 	           ?      # "   @ 	        3   A         1  	 B        7   C 	 	    % '   D  
         E +     *  +   F +     + C   G      " !   H &        &    I      0 .   J      ) (  
 K      ,    L      . /   M      4 5   N      6 5 ;   O  "    8 7 9   P  (    9 :   Q  $    < F   R 	 $       <   S +     > ?   T  $       =   U + .    ? @   V  .    @ A   W  *    A B   X      C , D   Y      D E   Z      F ; G   [ +     H  I   \ +     I J   ]      J K   ^      K L   _      L M   `      M N         3   Part 7 & 8  8  L   A* = a'bc' + a'b'c  8  L   B* = a'c' + a'b' + abc       C     Clock     PE     A     B                      P xd       �An                                                        