     
 LS Library                                   �          A                            
 LS Library                                  �        B                            
 LS Library                                  �        C                            
 LS Library          $                        �        D                            =
 LS Library         $                        �         ��         ��    �        ��      =
 LS Library                                 �         B�         B�    �        ��      =
 LS Library                                 �         b�         b�    �      	  ��      =
 LS Library                                  �         b�         b�    �   
     ��      D
 LS Library       ,                         �         ��         ��    �         ��         ��    �         ^         ^    �              ��      	 D
 LS Library       ,                         �         r�         r�    �         ��         ��    �   	      �         �    �              ��      
 M
 LS Library       9                         �   	      �3         �3    �   
      �1         �1    �           ��(       
 LS Library         @  
      ��         ��    �        e                                                                                    	         	         	                    
    	  	    
   
  
                                   
    	   
                          ! &  !   	 "  " #  #    $  $ %  %     &  &  ' '                                     	     %       
      %       
    % %                    	    %                        	 %           
               %            ,            ,           ,           1            ,   	         ,   	        ,   	        1   	       	  9   
         9   
      	  >   
        
  @           
  8          8          8        	  8        	  +          +                                & %        ! &         " *         # *         $ )         % )         & &                1   7-SEGMENT DISPLAY (e)        A      B     C     D     e                      P xd       �An                                                        