     
 LS Library	  	     -         ^I         ^I    �         3         3    �         �         �    �         .�         .�    �         b�         b�    �         ��         ��    �         \�         \�    �         �s         �s    �         �>         �>    �   	      �S         �S    �   
      �H         �H    �         jy         jy    �         >T         >T    �         Җ         Җ    �   A                           8  9  :  ;  <  �� |��C 4-BITFA.CKT C:\4-BITFA.CKT 4-BITFA.CKTa1  �V�    b1  �V�   a2  �V�   b2  �V�   a3  �V�   b3  �V�   a4  �V�  	 b4  �V�  
 C-in1 �V�   S1 n1 �V�    S2 n1 �V�   S3 n1 �V�   S4 n1 �V�   C-out4 V�   ���������������������������� �� �� �� ��
 ��	 �� �� �� �� �� �� �� �� ��    
 LS Library                6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                 �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �         ޗ         ޗ    �         t�         t�    �          ��         ��    �         �>         �>    �              	  �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �   	      ޗ         ޗ    �   
      t�         t�    �         ��         ��    �         �>         �>    �   
             �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library        "       6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ����������������������������                    ��        ��                   ��        ��       ��       ��        ��   	     ��  
     ��                 ��       ��       ��        ��       ��   
 LS Library         :  	      �]         �]    �         S1                            
 LS Library         :  
      ��         ��    �        S2                            
 LS Library         :        �         �    �        S3                            
 LS Library         :        �         �    �        S4                            
 LS Library         :        <�         <�    �        C-out                         
 LS Library                                  �        C-in                         
 LS Library                                  �        b1                           
 LS Library                                   �   @     a1                          	 
 LS Library                                  �        a2                          
 
 LS Library                                  �     	   b2                           
 LS Library                                  �      
   a3                           
 LS Library                                  �   !     b3                           
 LS Library                                  �   "     a4                           
 LS Library                                  �   #     b4                           ]
 LS Library                                �         "�         "�    �         �         �    �   ,   -   .  ��3        ]
 LS Library                                �         "�         "�    �         �         �    �   /   0   1  ��3        ]
 LS Library                                �         "�         "�    �         �         �    �   2   3   4  ��3        ]
 LS Library                                �         "�         "�    �         �         �    �   5   6   7  ��3                                     	                                                                                	           
                                                   
                         4 3   .      4   @ $  # 6   
   	     	  	 
  
       ! 3  <    0   -  ;   & ,  ' &  :   ' /  ( '  9   ( 2  ) (  8   ) 5  * &  + *  +    *        !  ? " ?  #   $ 1  %   &   '   = ( = > ) >  * % A + $ % ,   - "   . B   / B  0 7 C 1 D C 2 D  ��G E   +     - .    -             -        #    -        &    -        )    -        ,    -        /    -        2    -           	 7         
 8     	     9     
     7          )     % &    :          	  :          
  :        
    :        	    :            8          )     $ %    9          *     # "    :        
  *      ,    +            	           +                       *          '   	     !       
          '        '   !            " '        -   #            $ ,      +    % ,     * +    &           '           (           )          *  	         + - 	        ,            -           .             /            0           1         $   2            3           4            5            6           7         0   8 5           	 9 5          
 : 5           ; 5           < 5           = (     ' (   > (     ( )   ? *     ! "   @ '            A -         *    B +     . /   C ,     0 1   D ,     1 2   ����    "  6   4-bit Add/Subtract  
    " 1 - Subtract (A-B)
0 - Add (A+B)       S1     S2     S3     S4     C-out     C-in     b1     a1   	  a2 	 	 
  b2 
 
   a3     b3     a4     b4                                 	 	  
 
            P xd       �An                                                        