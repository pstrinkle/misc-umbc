      Generic Library                                 �         ~         ~    �         .         .    �         �         �    �         �         �    �      �@N W     �@N W   �      �@N W     �@N W   �                       ��   Generic Library                                   �         Asyn_Set                      Generic Library                                  �    
    FF_SET                        Generic Library          !                        �   	 
   Clk0                          �Bn        HBn       Clk0  Generic Library                                  �        FF_RESET                      Generic Library         &        r�         r�    �        Q                              Generic Library         &        ��         ��    �        QB                             Generic Library                                  �        Asyn_Reset                                                                                                     
     
                  	   
    	                                                                         	                                                                 	  "          
                                          	                              
     "    
     &            &            "          "          "          "                                          Asyn_Set     FF_SET     Clk0     FF_RESET     Q     QB    
 Asyn_Reset                            A �L       �An                                                         