     
 LS Library                                   �          A                            
 LS Library                                  �        B                            
 LS Library                                  �        C                            
 LS Library          $                        �        D                            =
 LS Library       $ $                        �         ��         ��    �        ��      =
 LS Library       $                         �         Ɛ         Ɛ    �        ��      =
 LS Library       $                         �         ��         ��    �      	  ��      =
 LS Library       $                          �         �T         �T    �   
     ��      D
 LS Library       0                         �         �         �    �         b�         b�    �         �         �    �              ��      	 D
 LS Library       0                         �         ��         ��    �         ��         ��    �   	      B�         B�    �              ��      
 D
 LS Library       0                         �         ��         ��    �         ^7         ^7    �   
      �"         �"    �              ��       D
 LS Library       0 $                        �         Z�         Z�    �          i         i    �         *g         *g    �              ��       M
 LS Library       8                         �   	      �j         �j    �         �         �    �   -   .   /  ��(       M
 LS Library       8   
                       �         �l         �l    �         �,         �,    �   0   1   2  ��(       M
 LS Library       @                         �         lC         lC    �         �~         �~    �   3   4   5  ��(       
 LS Library         H                         �   6     f                                                          
                             	   
            	                          	    
              	  	       
  
                                              . .     (                          	  " 
          !  !   "   "    $  # '  #   ! %  %    &  &   $ '  '   
 (  	 )  ( *  *   ) +  +    ,   ,  !  7 " 7 - # 8  $ 8 . %  9 & 9 0 ' :  ( : 1 ) ; 2 * ; 4 + / < , < 3 - 5 6 = =                                           %           $ %           ) %           $            )            $           	 )           
 $             )            0            0           0       
    5        !    0   	         0   	        0   	        5   	     #  	  0   
         0   
        0   
        5   
     %  
  0 %           0 &           0 '           5 &       '    "            "          -           -     	 
     /          ! /          " -     	     # ,         $ , %        % /         & "         ' ,          ( #            ) .         * # '         + . %        , - &         - 8        "   . 8       $  	 / =        +   0 8 !       &  
 1 8 #      (   2 = "       )   3 @        ,   4 @       *   5 E        -   6 H        -   7 5     ! "   8 5     # $  	 9 5 !    % &  
 : 5 #    ' (   ; =     ) *   < =     + ,         3   7-SEGMENT DISPLAY (f)        A      B     C     D     f                      P xd       �An                                                        