     
 LS Library                                   �          A                            
 LS Library                                  �        B                            
 LS Library                                   �        C                            
 LS Library          (                        �        D                            =
 LS Library                                  �         B�         B�    �        ��      =
 LS Library                                 �         B�         B�    �        ��      =
 LS Library                                  �         �T         �T    �      	  ��      =
 LS Library         (                        �         ��         ��    �   
     ��      A
 LS Library       ,                         �         Ɛ         Ɛ    �         r�         r�    �           ��      	 D
 LS Library       ,                         �         �         �    �         j�         j�    �   	      �3         �3    �              ��      
 D
 LS Library       ,                          �         �/         �/    �         "�         "�    �   
      Z�         Z�    �              ��       D
 LS Library       ,                          �         *g         *g    �         �          �     �         �j         �j    �              ��       M
 LS Library       4                         �         �l         �l    �         �j         �j    �   -   .   /  ��(       M
 LS Library       4  	                       �   
      �l         �l    �         �,         �,    �   0   1   2  ��(       M
 LS Library       =                         �         |r         |r    �         lC         lC    �   3   4   5  ��(       
 LS Library         C                         �   =     a                                                        	                          	             	             
             
         
            	  	        
  
                                              / /    '  , (  + )  !   
    "     $     	 % # 
 & %            !   "   #   $   %    '  	 (   )   &               *    *   )    +   (    ,  !  6 " 6 7 # 7 - $ 8  % 8 . &  9 ' 9 0 ( :  ) : 1 * ; 2 + ; 4 , / < - < 3 . 5 = > >                               !            )                         %                         %              !          	 % !          
   )           % )           ,            ,           1        $    ,   	         ,   	        ,   	        1   	     &  	  , !  
         , "  
        , #  
        1 "  
     (  
  ,             ,           ,            1        !     )                      !          ( #          ) "          * !        !          "          # +      	   $          % +      
 	   & +      
   ' ( )         ( ) !         ) *          *           + *         , )          - 4        #   . 4       %   / 9        ,   0 4        '  	 1 4       )  
 2 9        *   3 =        -   4 =       +   5 B        .   6 3     ! "   7 3     " #   8 1     $ %   9 1     & '  	 : 1     ( )  
 ; 9     * +   < 9     , -   = C        .       #  7 	  7-SEGMENT DISPLAY (a)        A      B     C     D     a                      P xd       �An                                                        