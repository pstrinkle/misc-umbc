 5 4   
 LS Library                                   �         C-in                         
 LS Library 	  	    ,        �@         �@    �         |/         |/    �         ,+         ,+    �         �t         �t    �         $         $    �         �         �    �         �         �    �         ��         ��    �   	      8         8    �   
      ��         ��    �         �          �     �         �"         �"    �         l*         l*    �         L(         L(    �         t�         t�    �          �-         �-    �         ��         ��    �         �         �    �         L         L    �         �         �    �         �         �    �         ��         ��    �         \         \    �         �         �    �         �         �    �         <         <    �                                                      
  	                �� ���C 8-BITFA.CKT C:\CIRCUITS\8-BITFA.CKT 8-BITFA.CKTa1  '�    b1  '�   a2  '�   b2  '�   a3  '�   b3  '�   a4  '�  	 b4  '�  
 b8  '�   a8  '�	   b7  '�
   a7  '�   b6  '�   a6  '�   b5  '�   C-in  '�   a5 n  '�   S1 n  '�    S2 n  '�   S3 n  '�   S4 n  '�   S5 n  '�   S6 n  '�   S7 n  '�   S8 n  '�  	 C-out '�  
 ����������������������������������������������������  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� ��    
 LS Library	  	     ! 	        ��         ��    �         �]         �]    �         lm         lm    �         m         m    �         
F         
F    �         ��         ��    �         b�         b�    �         ��         ��    �         �         �    �   	      �*         �*    �   
      &�         &�    �         ��         ��    �         F�         F�    �         
         
    �                               	  
        �� |��C 4-BITFA.CKT C:\4-BITFA.CKT 4-BITFA.CKTa1  �V�    b1  �V�   a2  �V�   b2  �V�   a3  �V�   b3  �V�   a4  �V�  	 b4  �V�  
 C-in1 �V�   S1 n1 �V�    S2 n1 �V�   S3 n1 �V�   S4 n1 �V�   C-out4 V�   ���������������������������� �� �� �� ��
 ��	 �� �� �� �� �� �� �� �� ��    
 LS Library                6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                 �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �         ޗ         ޗ    �         t�         t�    �          ��         ��    �         �>         �>    �              	  �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �   	      ޗ         ޗ    �   
      t�         t�    �         ��         ��    �         �>         �>    �   
             �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library        "       6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ����������������������������                    ��        ��                   ��        ��       ��       ��        ��   	     ��  
     ��                 ��       ��       ��        ��       ��  ���������������������������������������������������� 
 LS Library	  	     "        ��         ��    �         �]         �]    �         lm         lm    �         m         m    �         
F         
F    �         ��         ��    �         b�         b�    �         ��         ��    �         �         �    �         �*         �*    �         &�         &�    �         ��         ��    �         F�         F�    �         
         
    �   5   4   3   2   1   0   /   .                �� |��C 4-BITFA.CKT C:\4-BITFA.CKT 4-BITFA.CKTa1  �V�    b1  �V�   a2  �V�   b2  �V�   a3  �V�   b3  �V�   a4  �V�  	 b4  �V�  
 C-in1 �V�   S1 n1 �V�    S2 n1 �V�   S3 n1 �V�   S4 n1 �V�   C-out4 V�   ���������������������������� �� �� �� ��
 ��	 �� �� �� �� �� �� �� �� ��    
 LS Library                6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                 �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �         ޗ         ޗ    �         t�         t�    �          ��         ��    �         �>         �>    �              	  �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library               6�         6�    �   	      ޗ         ޗ    �   
      t�         t�    �         ��         ��    �         �>         �>    �   
             �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��    
 LS Library        "       6�         6�    �         ޗ         ޗ    �         t�         t�    �         ��         ��    �         �>         �>    �                �� ���C FA.CKT	 C:\FA.CKT FA.CKTC-in  �V�    Y in  �V�   X in  �V�   C-out �V�    Sum t �V�   ���������� �� ��  �� ��
 �� 	   :
 LS Library       $                          �         �,         �,    �         F,         F,    �            ��      :
 LS Library       $                         �         `�         `�    �         
A         
A    �           ��      :
 LS Library                                 �         �`         �`    �         �`         �`    �           ��     ������ :
 LS Library       ,                         �         �!         �!    �         j!         j!    �           ��      :
 LS Library       @                         �         �         �    �         r         r    �           ��      :
 LS Library       @                         �         ��         ��    �   	      :�         :�    �           ��     	 :
 LS Library       H                         �   	      ��         ��    �   
      ��         ��    �            ��     
 :
 LS Library       8                         �         &�         &�    �         ��         ��    �   !   "   #  ��      :
 LS Library       @                         �         l�         l�    �         �         �    �   /   0   1  ��     ����          ��                                       ��                ��      
             
         
                  	    	      	   
  	    ��        ��   ����������������������������                    ��        ��                   ��        ��       ��       ��        ��   	     ��  
     ��                 ��       ��       ��        ��       ��  ����          ��         ��        ��        ��        ��        ��        ��        ��        ��  	       ��   
      ��        ��        ��             ��       �� 	      �� 
      ��       ��       ��       ��           ��        ��       ��       ��       ��       ��   
 LS Library                                  �         A1                           
 LS Library                                  �        B1                           
 LS Library                                  �        A2                           
 LS Library                                  �        B2                           
 LS Library                                  �        A3                           
 LS Library                                  �         B3                           
 LS Library                                  �   !     A4                          	 
 LS Library                                  �   "     B4                          
 
 LS Library                                  �   #  	   A5                           
 LS Library                                  �   $  
   B5                           
 LS Library                                   �   %     A6                           
 LS Library                                  �   &     B6                           
 LS Library          $                        �   '     A7                           
 LS Library          #                         �   (     B7                           
 LS Library          ( 
                       �   )     A8                           
 LS Library          ' !                       �   *     B8                           
 LS Library         ;        ��         ��    �   +     S1                            
 LS Library         ;        ��         ��    �   ,     S2                            
 LS Library         ;         �          �    �   -     S3                            
 LS Library         ;        Z�         Z�    �   .     S4                            
 LS Library         ;        ��         ��    �   /     S5                            
 LS Library         ;        ��         ��    �   0     S6                            
 LS Library         ;        �         �    �   1     S7                            
 LS Library         ;        B�         B�    �   2     S8                            ]
 LS Library        	                         �         dR         dR    �         ��         ��    �   B   C   D  ��3        
 LS Library         8         ��         ��    �   4     C-out                         ]
 LS Library                                 �         B	         B	    �         ��         ��    �   E   F   G  ��3        ]
 LS Library                                 �         ��         ��    �         ��         ��    �   H   I   J  ��3        ]
 LS Library                                 �         "�         "�    �         J         J    �   K   L   M  ��3        ]
 LS Library                                 �         �         �    �         �
         �
    �   N   O   P  ��3         ]
 LS Library                                 �         |t         |t    �         ��         ��    �   Q   R   S  ��3       ! ]
 LS Library        !                         �          ��         ��    �         L�         L�    �   T   U   V  ��3       " ]
 LS Library        %                         �   !      �o         �o    �   	      ��         ��    �   W   X   Y  ��3       # 
 LS Library	  	     $ 4 "                       �   #      n;         n;    �   $      ;         ;    �   %      �:         �:    �   &      ~:         ~:    �   '      .:         .:    �   (      �9         �9    �   )      �9         �9    �   *      >9         >9    �   +     N �8        N �8    �   ,      �8         �8    �   -      N8         N8    �   .      �7         �7    �   /      �7         �7    �   �   �   �   �   �   �   �   �   �   �  �  �  �  �  ��1 $ 
 LS Library          5 "                       �   #      
         
    �   $      �         �    �   %      j         j    �   0                   �   1      �         �    �   2      z         z    �   3      *         *    �   �    X                           % 
 LS Library          : 4                       �   5      F�         F�    �   6      ��         ��    �   7      ��         ��    �   8      V�         V�    �   9      �         �    �   :      ��         ��    �   ;      f�         f�    �   �    Y                           & 
 LS Library          7 *      \�         \�    �   �     Cin                         ' `
 LS Library       6 "      ~         ~    �   #      $         $    �   $      �,         �,    �   %      �M         �M    �   0      ZV         ZV    �   1      �^         �^    �   2      ~g         ~g    �   3       r          r    �   "      �|         �|    �   #      ��         ��    �   $      �I         �I    �   %      Z�         Z�    �   0      ��         ��    �   1                   �   2      �          �     �   3      &)         &)    �   �  �  �   ��                                               ( `
 LS Library       : &      �G         �G    �   '      �G         �G    �   (      �S         �S    �   )      ZS         ZS    �   <      
S         
S    �   =      �R         �R    �   >      ]         ]    �   ?      �\         �\    �   &      h\         h\    �   '      \         \    �   (      �[         �[    �   )      x[         x[    �   <      ([         ([    �   =      �e         �e    �   >      Je         Je    �   ?      �d         �d    �   �  �  �   ��                                               ��* `
 LS Library      ! 6 "      �c         �c    �   #      �m         �m    �   $      hm         hm    �   %      m         m    �   "      �l         �l    �   #      xl         xl    �   $      (l         (l    �   %      �k         �k    �   �  �  �  �  �   ��
                                            + `
 LS Library      ! : &      �z         �z    �   '      Nz         Nz    �   (      �y         �y    �   )      �y         �y    �   &      ^y         ^y    �   '      y         y    �   (      �x         �x    �   )      nx         nx    �   �  �  �  �  �   ��
                                            , `
 LS Library       * 8 +      x         x    �   ,      �w         �w    �   -      ~w         ~w    �   .      .w         .w    �   +      �v         �v    �   ,      �v         �v    �   -      >v         >v    �   .      ��         ��    �   �   �   �   �   �  ��                                            - 
 LS Library	        8 4      Z�         Z�    �   5      tb         tb    �   6      �a         �a    �   7      4a         4a    �   8      �`         �`    �   9      �_         �_    �   :      T_         T_    �   ;      �^         �^    �   *      �R         �R    �   &      J         J    �   '      4I         4I    �   (      �O         �O    �   )      �N         �N    �   <      ^N         ^N    �   =      �M         �M    �   >      �]         �]    �   ?      $]         $]    �   �   �   �  �� 6��C 8-BITXOR.CKT C:\CIRCUITS\8-BITXOR.CKT 8-BITXOR.CKTB �</�</    C-in �</   XOR'd �</    ����������������������������������  �� �� �� �� �� �� �� �� ��	 ��
 �� �� �� �� �� �� �� 
 ���� ]
 LS Library                                  �         t�         t�    �   	      $�         $�    �           ��3        ]
 LS Library                                 �         ��         ��    �   
      ��         ��    �           ��3        ]
 LS Library                                 �         D�         D�    �         �         �    �      	   
  ��3        ]
 LS Library         %                        �         �y         �y    �         By         By    �           ��3        ]
 LS Library         +                        �         �k         �k    �         �k         �k    �           ��3        ]
 LS Library         0                        �         .^         .^    �         �]         �]    �           ��3        ]
 LS Library         6                        �         |P         |P    �         ,P         ,P    �           ��3       	 ]
 LS Library         ;                        �         �B         �B    �         zB         zB    �           ��3       
 `
 LS Library               8�         8�    �         �         �    �         �I         �I    �         �I         �I    �         >I         >I    �         �H         �H    �         �H         �H    �         NH         NH    �          �G         �G    �         �G         �G    �         ^G         ^G    �         G         G    �         �F         �F    �         nF         nF    �         F         F    �         �E         �E    �                  !      ��                                                                                 `
 LS Library       0  	      �D         �D    �   
      �B         �B    �         ~B         ~B    �         .B         .B    �         �A         �A    �         �A         �A    �         >A         >A    �         �@         �@    �   	      �@         �@    �   
      N@         N@    �         �?         �?    �         �?         �?    �         ^?         ^?    �         ?         ?    �         �>         �>    �         n>         n>    �   9   :   ;   <   =   >   ?   @   A  ��                                                                                ��     ��         ��        ��        ��        ��        ��        ��        ��  	     	 ��                       	   	      ��   
      ��        ��        ��        ��        ��        ��    	    ��  . `
 LS Library       > 3 +      ��         ��    �   ,      v�         v�    �   -      &�         &�    �   .      ��         ��    �   @      ��         ��    �   A      6�         6�    �   B      ��         ��    �   C      ��         ��    �   +      ��         ��    �   ,      ��         ��    �   -      Z�         Z�    �   .      
�         
�    �   @      ��         ��    �   A      j�         j�    �   B      �         �    �   C      ��         ��    �   �   �   �  ��                                               / 
 LS Library         = < D      �C         �C    �   �     Cout                         0 
 LS Library         A 2 +      �>         �>    �   ,      �<         �<    �   -      �<         �<    �   .      F<         F<    �   @      �;         �;    �   A      �;         �;    �   B      V;         V;    �   C      ;         ;    �   �     Sum                          1 
 LS Library	  	     2 5 0                       �   1      n;         n;    �   2      ;         ;    �   3      �:         �:    �   <      ~:         ~:    �   =      .:         .:    �   >      �9         �9    �   ?      �9         �9    �   /      >9         >9    �   @     N �8        N �8    �   A      �8         �8    �   B      N8         N8    �   C      �7         �7    �   D      �7         �7    �   �   �   �   �   �   �   �   �   �   �  �  �  �  �  ��1 2 `
 LS Library      / ; <      F�         F�    �   =      ��         ��    �   >      ��         ��    �   ?      V�         V�    �   <      �         �    �   =      ��         ��    �   >      f�         f�    �   ?      �         �    �   �  �  �  �  �   ��
                                            3 `
 LS Library      / 7 0      ��         ��    �   1      v�         v�    �   2      &�         &�    �   3      ��         ��    �   0      ��         ��    �   1      6�         6�    �   2      ��         ��    �   3      ��         ��    �   �  �  �  �  �   ��
                                            4 `
 LS Library       8 9 @      F�         F�    �   A      ��         ��    �   B      ��         ��    �   C      V�         V�    �   @      �         �    �   A      ��         ��    �   B      f�         f�    �   C      �         �    �   �   �   �   �   �  ��                                            E E   
         "    !                                                                                                      	     "    
    	         
 !                                              
                                                                                                                   	                                 !   !      "   "  #    $    #  #   $   $  #   $   %  #   $   &  #   -    '  #   -   (  #   -   )  #   -   *  #   -   &    +  #    0    ,  #   0   -  #   0   .  #   0   /  #   1   0  $   1    1  $   1   2  $   1   3  $   1   4  %    -    5  %   -   6  %   -   7  %   -   8  %   -   9  %   -   :  %   -   ;  %   -   <  -   1   =  -   1   >  -   1   ?  -   1   @  1    0   A  1   0   B  1   0   C  1   0   D  1   /    ~ ~   
 +  3 /  5 3   5  6 .  7 6   7  8 -  9 8 	  9 
 : ,  	 :   ;  ; <  < 0   =  = >  > 1   ?  ? @  @ 2   A  A 4  \ [  \ W  ] c  ^ ]  ^    ]  [ T  [ Z  Z Q   Z _ ! _ N " _ ` # ` K $ ` a % a H & a b ' b E ( b c ) c B *  F +  C ,   I - $ O . " L / & R 0 ( U 1 * X 2 e  3 e f 4 S f 5 g  6 g h 7 % h 8 i  9 i j : P j ; k  < k l = # l > m  ? m n @ M n A o  B p o C q p D q r E ! r F s  G t s H J t I u  J v u K w v L w  M y  N x y O   P G x Q z  R { z S D { T |  U } | V   } W ' d X ~ d Y ~  Z V  [ �  \ �  ] ) � ^ � � _ �  ` Y � a � � b �  c � � d � � e � � f � � g � � h � � i � � j � � k � � l � � m � � n � � o � � p � � q � � r � � s � � t � � u � � v � � w � � x � � y � � z � � { � � | � � } � � � �           V                  4           4           4           4           4           4           4       	   	 4          
 4             ,       ;    ,            ,       8    ,       5    ,       2    ,       Y    ,     
  \    ,     	  _  
  ,       b  	  ,       >    ,       A    ,       F    ,       I    ,       M    ,       O    ,       Q    ,        T            +            O            *            L             ,   !         E   "    	     .   #    
     =   $         -   %  !       7   &          /   '  %       W   (  $       0    )  )       ]  
 *  (       1  ! + ;            , ;        
   - ;           . ;           / ;           0 ;           1 ;           2 ;           3 8         4 8 !          5 8         6 9         7 9         8 :         9 :     	    : ;      
   ; 7         < 7         = 6         > 6         ? 5         @ 5         A 4 !        B  
       )    C        +   D         S   E         '    F        *   G         P   H         %    I        ,   J         H   K         #    L        .   M         @   N         !    O        -   P         :   Q              R          /   S          4   T  "  !         U  $  !    0    V  #  !     Z   W  &  "         X  (  "    1  ! Y  '  "     `  	 Z             [  "          \  &         ]            ^ ,          _        ! "    `      " # $    a      $ % &    b      & ' (    c  
    (  )    d % %    W X   e $     3 2   f $     4 3   g #     6 5   h # !    7 6   i "     9 8   j "     : 9   k !     < ;   l !     = <   m       ? >   n       @ ?   o &     B A   p &     C B   q      D C   r      E D   s '     G F   t '     H G   u (     J I   v (     K J   w      L K   x )     P N   y )     N M   z *     R Q   { *     S R   | +     U T   } +     V U   ~ %     X Y    & #    Z [   � &     [ \   � ' )    ] ^  
 � '     ^ _  
 � ( '    ` a  	 � (     a b  	 � $ 6  #    *       " � $ 7  #   *      # � $ 8  #   *      $ � $ 9  #   *      % � $ :  #   +       & � $ ;  #   +      ' � $ <  #   +      ( � $ =  #   +      ) � $ >  #    }  * � * 8  #    ,       + � * 9  #   ,      , � * :  #   ,      - � * ;  #   ,      . � * <  #    {  / �  6  $     z  " # $ % 0 1 2 3 �  ;  %     f  4 5 6 7 8 9 : ; �  8  &     e  * �  6  '     y  " # $ % �  7  '    x  0 1 2 3 �  :  (     w  & ' ( ) �  ;  (    v  < = > ? �����  >    | }  * �  8    c e |  * �  6  '     z  " # $ % 0 1 2 3 �  :  -    (       & ' ( ) < = > ? �  :  -    d  * �  8    d c  * �  ;  -     f  4 5 6 7 8 9 : ; � ! 6  *     y  " # $ % � ! :  +     w  & ' ( ) � - 8  ,     u  + , - . � ; 4    h g  @ A B C � . 3    j i  + , - . � 2 7  1    3       0 � 2 8  1   3      1 � 2 9  1   3      2 � 2 :  1   3      3 � 2 ;  1   2       < � 2 <  1   2      = � 2 =  1   2      > � 2 >  1   2      ? � 2 ?  1    q  / � 8 9  1    4       @ � 8 :  1   4      A � 8 ;  1   4      B � 8 <  1   4      C � 8 =  1    p  D �   2    l k  0 1 2 3 � - 7    n m  0 1 2 3 � - 2    n l  0 1 2 3 �   @    r o  < = > ? � / ;  2     s  < = > ? � - @    t r  < = > ? � - ;    t s  < = > ? � . 8    u j  + , - . �   ;    v o  < = > ? �   7    x k  0 1 2 3 � A 3  .    0       + , - . @ A B C � / 7  3     m  0 1 2 3 � > 4  .    h  @ A B C � > 3  .     i  + , - . � ; 9  4     g  @ A B C � = =  /     p  D � * ?    { q  /     (  <   8-Bit Full Adder/Subtractor      + Part 1: 
8th Bit is more Significant(128)   0  2  Part 2         C-in      A1     B1     A2     B2     A3     B3     A4   	  B4 	 	 
  A5 
 
   B5     A6     B6     A7     B7     A8     B8     S1     S2     S3     S4     S5     S6     S7     S8   $  X $    C-out   %  Y %  &  Cin & �� /  Cout /  0  Sum 0                                	 	  
 
                                                               P xd      �An                                                        