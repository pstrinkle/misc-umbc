     u            u Generic Library       )                           �         6�         6�    �         R�         R�    �         �         �    �         ��         ��    �         D�         D�    �        +       
  ��      �AN        �@N          Meg         �<N1  Generic Library          (                        �   ) 
    Clk0                          �Bn        HBn       Clk0 u           u Generic Library       (                          �         ��         ��    �         ��         ��    �         $�         $�    �         l�         l�    �         ��         ��    �   2     *         ��      �AN        �@N          Meg         �<N1  Generic Library           	                       �   	     C                            A Generic Library       #                         �   
      ��         ��    �         ��         ��    �   !         ��-       ] Generic Library         	                       �         F�         F�    �   
      v�         v�    �   3   1   0  ��M        ] Generic Library       "                          �         ��         ��    �         ��         ��    �      $   %  ��M        A Generic Library        !                        �   	      ��         ��    �         ��         ��    �   &   '   (  ��-        Generic Library         4         t          t    �        A                            	  Generic Library         4 !       Zo         Zo    �   ,     B                            
  Generic Library                                   �    
    SetHigh                       Generic Library          
                        �        SetHigh2                                  
                                                      	                                          	             
                  * *                      +       	   
  !              0    " 3  " #  ' #  / 1  	      %   )    .     ( $  /    ,   -  - #      . & ! *  " 2  #   $    %    &  4 ' 4  ( 4 5 ) 5  6 6   /      $ %     0 "          /     # $     +     "   #     + 	                   &    4             	  
          ! !        	           	 
 / #           / "            , &       )    !          ) "           ,          %     ( #     !     .           1          (               ( )         .        	    +       '    1     	      0                  	  " !                      !      
    !          0          0           #         
 ! #        
   "         	 #  $        	 $ " #         % ' "          &  "           '  $        	 ( ! #          )  )          * (       !   + ) #          , 4 "  	        -  $       	 .  "         /          0 !          
 1           2 +        "    3           	 4      ' & (   5  &    ( )             Clk0     C     A   	  B 	  
  SetHigh 
    SetHigh2                         P xd       �An                                                        