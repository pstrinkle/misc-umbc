     
 LS Library          $                         �          D                            
 LS Library                                  �        C                            
 LS Library                                  �        B                            
 LS Library                                  �        A                            =
 LS Library        $                         �         �,         �,    �        ��      =
 LS Library                                �         �j         �j    �        ��     �� =
 LS Library                                �         �j         �j    �   
     ��      =
 LS Library                                �         *g         *g    �        ��     	 A
 LS Library       (                         �         Z�         Z�    �         "�         "�    �           ��      
 A
 LS Library       (                         �          �1         �1    �   	      �3         �3    �           ��       D
 LS Library       (                         �         �         �    �         ��         ��    �   
      r�         r�    �              ��       D
 LS Library       ( $                        �         ^         ^    �         ��         ��    �         ��         ��    �              ��       M
 LS Library       0   
                       �         b�         b�    �         �         �    �           ��(       M
 LS Library       0                         �   	      �         �    �         B�         B�    �          !  ��(       M
 LS Library       8                         �         ��         ��    �         B�         B�    �   "   #   $  ��(       
 LS Library         ?                         �   F     c                                          
                       	                                                         	    
      	        	  
       
                                                6 6       &   =    )   (  
 &  % &  %   B A 	 + B 
 *    )  * )   ,  -   . -   .   .  ( '  '    /  0 /  0   ! 2  2 1  1 "   3  4 3  4 #   5  6 5  6      7 ! 7 8 " 8  #  9 $ 9 : % :  &  ; ' < ; ( <  )  = * = > + > ? , @ ? - @  . , + /  B 0 A  1 ' C 2 C D 3 E D 4 E  5 $ F G E    %                                                   %            ! %                        !           ����
             !                    )    !            (   	         (   	        -   	          (   
         (   
    
     -   
       	  (        /    (           (           -        #  
  ( %       -    ( &      0    ( '      4    - &       &    0 !       %  
  0 #      (    5 "           0        "     0         	 ! 5           " 8           # 8          $ =        5   %          &           ' %       1   ( %         )  %          *       
    + &     . 	   , &      .   - '         . '          / $ %        0 $         1 7         2 7         3 7 "        4 7         5 /        	 6 /        	 7 /       !   8 /     ! "   9 /     # $  
 : / !    $ %  
 ; / &    & '   < / #    ' (   =      )  *   >  '    * +   ? & '    + ,   @ & %    , -   A ' &     0   B '     / 	    C % (    1 2   D ' (    2 3   E ' '    3 4   F ?        5         2   7-SEGMENT DISPLAY (c)        D      C     B     A     c                      P xd       �An                                                        